--------------------------------------------------------------------------------
-- Energy Detection UWB Receiver TESTBENCH  
-- PSBC Final project A.A. 2007-2008  
--
-- Testbench which generates input signals and the expected outputs
-- for the digital backend/memory encoder and decoder subsystems. 
-- 
-- "system" components is your final project including everything
-- memory, bus encoding/decoding, backend...  
--
-- Once simulation is run, the architecture creates the two files 
-- DATAIN.DAT and DATAOUT.DAT
-- 
-- The DATAIN.DAT file is generated by the testbench only and 
-- contains the correct data sequence which the digital system 
-- must produce...
--
-- The DATAOUT.DAT file includes the demodulated data given by
-- system component instantiation....
--
-- If DATAOUT.DAT and DATAIN.DAT match for a large number 
-- of clock cycles, your system is working correctly (with good probability)...
--------------------------------------------------------------------------------



-- IMPORTANT!!
-----------------------------------------------------------------
--
-- Guidelines for writing VHDL human readable code:
--
-- One of the most important aspects of hardware description
-- languages such as VHDL is the code portability. A good VHDL 
-- code is also a readlable and understandable. Follow these tips 
-- while creating each VHDL file:
--
-- USE AN ENTITY NAME SIMILAR TO THE SIGNAL OPERATION 
--   If you call the output enable signal "STAR" it will be 
--   very difficult for a new reader to understand...
-- COMMENT THE CODE
--   If between a modification to another you wait a long time, 
--   you will spend to much time re-understanding what the architecture
--   do... 
-- ADD A REVISION TABLE AT THE BEGINNING OF EACH VHDL FILE
--   Good VHDL files also have a "comment table" which includes e.g. 
--   the last modification date, the authors, the revision number, 
--   a brief description of the architecture and entity, and so on...
--   E.g.
--  -----------------------------------------
--   -- Authors: Behzad Razavi
--   -- Last modification: 02/10/2004
--   -- Revision: 1.3
--   -- Desc: High school project
--   --
--   -- Viterbi encoder, decodes SI input into
--   -- SO output using the Viterbi algorithms...
--   -- CLK = clock
--   -- RESET = reset
--   -- DIN = Data in (10 bits)... 
--   -- DOUT = Data out (Nb bits, see package 'definitions')
--  -----------------------------------------
--
--  -------------------------------------------
--   -- Authors: Colonna Alessandro, Cutrupi Massimo
--   -- Last modification: 11/03/2008
--   -- Revision: 1.0
--   -- Desc: Low-Power System Design project
--   --
--   -- UWB baseband processing power optimization
--   -- Digital-Backend + Bus Encoder/Decoder + Memory Multi-Banks & Multi-
--   -- Symbol for word optimization (see constants_def.vhd & array_def.vhd for
--   -- information)
--   --
--  -----------------------------------------
--
-- Whatever you want to add...
--
-----------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use ieee.math_real.all;  -- This is to use real signals... 
use ieee.numeric_std.all;
use std.textio.all;      -- This is to include the function for 
                         -- reading and writing files (e.g. dataout.dat)...
use ieee.std_logic_textio.all;
use work.constants_def.all;
-- use work.array_def.all;

-- A testbench has got any connection to the extern world... 
entity tb_system is
  
end tb_system;


-- it has only an architecture... 
architecture test of tb_system is

-- This is YOUR system component declaration... 
-- MAKE SURE your entity has the same names 
-- reported here... 

component UWB_system

  generic (
    M    : integer ;
    N    : integer ;
    NQ   : integer ;
    logM : integer ;
    logN : integer );

  port (
    ck_slow      : in  std_logic;
    ck           : in  std_logic;
    reset        : in  std_logic;
    start        : in  std_logic;
    DIN          : in  std_logic_vector(NQ-1 downto 0);
    DOUT         : out std_logic_vector(M-1 downto 0);
    DBUS         : out std_logic_vector(M-1 downto 0);
    MEMADDBUS    : out arr_add;
    MEMDATABUS   : out arr_data;
    GCLK_mem     : out std_logic_vector(NBANKS-1 downto 0);    
    voutset      : out std_logic);
    
end component;

component memory
  generic( DBITS: integer;             
           ABITS: integer);           
           --WORDS: integer:=1024);                         -- WORDS=2**ABITS

  port( DIN     : in  std_logic_vector(DBITS-1 downto 0); 	-- input data
        DOUT    : out std_logic_vector(DBITS-1 downto 0);       -- output data
        ADD     : in  std_logic_vector(ABITS-1 downto 0);  	-- addresses
	ck      : in  std_logic;
	WR      : in  std_logic;
        OE      : in  std_logic);
end component;


  signal int_DIN, int_DOUT: arr_data;
  signal int_ADD : arr_add;
  signal int_GCLK_mem : std_logic_vector(NBANKS-1 downto 0);

  signal ck : std_logic := '1';
  signal ck_slow: std_logic := '0';
  signal reset : std_logic := '0';
  signal start : std_logic := '0';

  signal voutset : std_logic := '0';
  constant NQ : integer := NQ;
  constant N : integer := N;
  constant M : integer := M;
  -- constant ABITS : integer := 2;
  signal DIN : std_logic_vector(NQ-1 downto 0) := (others => '1');
  signal DOUT : std_logic_vector(M-1 downto 0);
  signal DBUS : std_logic_vector(M-1 downto 0);

begin  -- test

 
  ck <= not ck after 0.5 ns;

  ck_slow_p: process (ck, reset)
  begin  -- process ck_slow_p
    if reset = '0' then                 -- asynchronous reset (active low)
      ck_slow<='0';
    elsif ck'event and ck = '1' then    -- rising clock edge
      if start='1' then
        ck_slow<=not(ck_slow);
      end if;
    end if;
  end process ck_slow_p;

  -- asynch reset
  reset <= '1', '0' after 0.1 ns, '1' after 0.2 ns; 

  -- start signal
  start <= '1' after 8.25 ns;
  
  -- DIN assignment
  pdin: process(ck,reset)
  variable ncntr,mcntr: integer :=0;
  variable seed1 : positive := 3565;
  variable seed2 : positive := 4523;
  variable awgn,x1,z1,z2 : real := 0.0;
  variable y1,z3 : integer := 0;
  constant sigma : real := 0.4;         -- awgn variance
  file datain : text is out "datain.dat";  -- input data
  variable fileline : line;
  begin
    if reset='0' then
      DIN <= (others => '0');
    elsif ck'event and ck='1' then
      if start='1' then
        if ncntr=0 then
          uniform(seed1,seed2,x1);  
          y1:=integer(trunc(x1*real(M)));
          write(fileline,y1);
          writeline(datain,fileline);
        end if;
        uniform(seed1,seed2,z1);        
        uniform(seed1,seed2,z2);
        awgn:=sigma*sqrt(-2.0*log(z1))*cos(2.0*math_pi*z2);
        if mcntr=y1 then
          z3:=integer(trunc((awgn+0.75*real(2**(NQ)))));
          -- saturation
          if z3>2**(NQ-1) then
            z3:=2**(NQ-1);
          end if;
          if z3<0 then
            z3:=0;
          end if;
          DIN <= std_logic_vector(to_unsigned(z3,DIN'length));
          -- DIN(0) <= '1';
        else
          z3:=integer(trunc(awgn));
          -- saturation
          if z3>2**(NQ-1) then
            z3:=2**(NQ-1);
          end if;
          if z3<0 then
            z3:=0;
          end if;         
          DIN <= std_logic_vector(to_unsigned(z3,DIN'length));
          -- DIN(0) <= '0';
        end if;
        mcntr:=(mcntr+1) mod M;
        ncntr:=(ncntr+1) mod (M*N);
      end if;
    end if;
  end process;

  -- DOUT output file
  -- Creates the output file reading information
  -- from DOUT...
  -- Make sure that your system includes the 'voutset' output signal...   
  pdout: process(ck)
  file dataout : text is out "dataout.dat";  -- output data
  variable fileline : line;
  begin
    if ck'event and ck='1' then
      if (voutset)='1' then
        for i in M-1 downto 0 loop
          if DOUT(i)='1' then
            write(fileline,i);
            writeline(dataout,fileline);
          end if;
        end loop;  -- i
      end if;
    end if;
  end process;
  
-- System instantiation... 
  system_inst: UWB_system
    generic map (
      N     => N,
      M     => M,
      NQ    => NQ,
      logM  => logM,
      logN  => logN)
    port map (
      ck_slow    => ck_slow,
      ck         => ck,      
      reset      => reset,
      start      => start,
      DIN        => DIN,
      DOUT       => DOUT,
      DBUS       => DBUS,
      MEMADDBUS  => int_ADD,
      MEMDATABUS => int_DIN,
      GCLK_mem   => int_GCLK_mem,   
      voutset    => voutset);

-- Memory instantiation... 
  mem_inst: for i in NBANKS-1 downto 0 generate
    inst_mem_banks : memory generic map (
      DBITS => NBIT1WORD,
      ABITS => NADD1BANK)
      port map (
        DIN 		=> int_DIN(i),
        DOUT            => int_DOUT(i),
        ADD             => int_ADD(i),
        ck              => int_GCLK_mem(i),
        WR              => '1',
        OE              => '1');
  end generate mem_inst;
   
end test;
